module basic_mux_tb();
   

   
endmodule